module Compare_Hash(
//	 input Clk, Reset,
 //   input reg[127:0]hash_in,
//	 output Result
);


endmodule
